20002.5